return {
-- Table: {1}
{
   ["soundVolume"]=0.01,
   ["fullScreen"]=false,
   ["uiZoomToggle"]=false,
},
}